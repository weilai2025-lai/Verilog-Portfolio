library verilog;
use verilog.vl_types.all;
entity accumulator_vlg_vec_tst is
end accumulator_vlg_vec_tst;
