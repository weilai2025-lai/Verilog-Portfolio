library verilog;
use verilog.vl_types.all;
entity fp_addfull_vlg_vec_tst is
end fp_addfull_vlg_vec_tst;
