library verilog;
use verilog.vl_types.all;
entity seven_seg_10_vlg_vec_tst is
end seven_seg_10_vlg_vec_tst;
