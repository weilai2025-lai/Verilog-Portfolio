library verilog;
use verilog.vl_types.all;
entity mem1_vlg_vec_tst is
end mem1_vlg_vec_tst;
