library verilog;
use verilog.vl_types.all;
entity count111_moore_vlg_vec_tst is
end count111_moore_vlg_vec_tst;
