library verilog;
use verilog.vl_types.all;
entity add6_vlg_vec_tst is
end add6_vlg_vec_tst;
