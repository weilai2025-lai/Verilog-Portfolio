library verilog;
use verilog.vl_types.all;
entity count111_improved_vlg_vec_tst is
end count111_improved_vlg_vec_tst;
