library verilog;
use verilog.vl_types.all;
entity mux8to1_vlg_vec_tst is
end mux8to1_vlg_vec_tst;
