library verilog;
use verilog.vl_types.all;
entity srdisplay_vlg_vec_tst is
end srdisplay_vlg_vec_tst;
