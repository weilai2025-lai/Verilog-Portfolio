library verilog;
use verilog.vl_types.all;
entity register_vlg_vec_tst is
end register_vlg_vec_tst;
