library verilog;
use verilog.vl_types.all;
entity D_Latch_vlg_vec_tst is
end D_Latch_vlg_vec_tst;
