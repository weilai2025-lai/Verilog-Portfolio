library verilog;
use verilog.vl_types.all;
entity SR_Latch_vlg_vec_tst is
end SR_Latch_vlg_vec_tst;
