library verilog;
use verilog.vl_types.all;
entity ffulladd_clg_vlg_vec_tst is
end ffulladd_clg_vlg_vec_tst;
