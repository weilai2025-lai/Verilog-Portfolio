library verilog;
use verilog.vl_types.all;
entity pencoder_8bit_vlg_vec_tst is
end pencoder_8bit_vlg_vec_tst;
