library verilog;
use verilog.vl_types.all;
entity seven_segnent_vlg_vec_tst is
end seven_segnent_vlg_vec_tst;
