library verilog;
use verilog.vl_types.all;
entity fulladd32bit_vlg_vec_tst is
end fulladd32bit_vlg_vec_tst;
