library verilog;
use verilog.vl_types.all;
entity SR_Latchbev_vlg_vec_tst is
end SR_Latchbev_vlg_vec_tst;
