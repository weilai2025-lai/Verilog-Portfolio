library verilog;
use verilog.vl_types.all;
entity fulladd16bit_vlg_vec_tst is
end fulladd16bit_vlg_vec_tst;
