library verilog;
use verilog.vl_types.all;
entity traffic_moore_vlg_vec_tst is
end traffic_moore_vlg_vec_tst;
