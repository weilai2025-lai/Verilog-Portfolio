library verilog;
use verilog.vl_types.all;
entity pencoder_4bit_vlg_vec_tst is
end pencoder_4bit_vlg_vec_tst;
