library verilog;
use verilog.vl_types.all;
entity ffulladd_cla_vlg_vec_tst is
end ffulladd_cla_vlg_vec_tst;
