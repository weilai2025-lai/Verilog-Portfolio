library verilog;
use verilog.vl_types.all;
entity AccumDC_vlg_vec_tst is
end AccumDC_vlg_vec_tst;
