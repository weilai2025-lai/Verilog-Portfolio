library verilog;
use verilog.vl_types.all;
entity traffic_moore2_vlg_vec_tst is
end traffic_moore2_vlg_vec_tst;
