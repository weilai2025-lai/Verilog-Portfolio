library verilog;
use verilog.vl_types.all;
entity stack_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        data_in         : in     vl_logic_vector(3 downto 0);
        enable          : in     vl_logic;
        push_pop        : in     vl_logic;
        rst             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end stack_vlg_sample_tst;
