library verilog;
use verilog.vl_types.all;
entity Dff_behavioral_vlg_vec_tst is
end Dff_behavioral_vlg_vec_tst;
