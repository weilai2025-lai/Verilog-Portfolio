library verilog;
use verilog.vl_types.all;
entity queue_vlg_vec_tst is
end queue_vlg_vec_tst;
