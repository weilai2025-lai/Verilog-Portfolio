module fulladd(a,b,cin,s,cout);
input a,b,cin;
output s,cout;

assign {cout,s}=a+b+cin;

endmodule

