library verilog;
use verilog.vl_types.all;
entity shiftreg_vlg_vec_tst is
end shiftreg_vlg_vec_tst;
