library verilog;
use verilog.vl_types.all;
entity div_decoder_vlg_vec_tst is
end div_decoder_vlg_vec_tst;
