library verilog;
use verilog.vl_types.all;
entity floating_adder_withsubtraction_vlg_vec_tst is
end floating_adder_withsubtraction_vlg_vec_tst;
