library verilog;
use verilog.vl_types.all;
entity Priority_encoder_vlg_vec_tst is
end Priority_encoder_vlg_vec_tst;
