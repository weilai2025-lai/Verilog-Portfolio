module div_dec(din, dout);

input [2:0]din;
output reg[31:0]dout;

always @(din)
begin
	case(din)
	3'd0: dout=32'd200000000;
	3'd1: dout=32'd150000000;
	3'd2: dout=32'd100000000;
	3'd3: dout=32'd50000000;
	3'd4: dout=32'd25000000;
	3'd5: dout=32'd166700000;
	3'd6: dout=32'd10000000;
	3'd7: dout=32'd4;
	endcase
end
endmodule

	
	