library verilog;
use verilog.vl_types.all;
entity FP_ADD_vlg_vec_tst is
end FP_ADD_vlg_vec_tst;
