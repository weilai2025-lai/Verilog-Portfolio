library verilog;
use verilog.vl_types.all;
entity fulladd_bev_vlg_vec_tst is
end fulladd_bev_vlg_vec_tst;
