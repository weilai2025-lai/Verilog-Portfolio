library verilog;
use verilog.vl_types.all;
entity stack_vlg_vec_tst is
end stack_vlg_vec_tst;
