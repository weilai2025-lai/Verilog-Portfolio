library verilog;
use verilog.vl_types.all;
entity bounce_avoid_vlg_vec_tst is
end bounce_avoid_vlg_vec_tst;
