module fp_addfull(fa,fb,fs,op);
parameter width_total = 32;
parameter width_e = 8;
parameter width_f = 23;

input op;
input [width_total-1:0]fa,fb;
output [width_total-1:0]fs;
wire valid,zero;
wire fa_s,fb_s,fs_s;
wire [width_total-1:0]fb_math;
wire [width_e-1:0]fa_e,fb_e,fs_e,ex_diff;
wire [width_f-1:0]fa_f,fb_f,fs_f;
wire [width_f+3-1:0]fa_fex,fb_fex,fs_fcal,fb_fexshift;
wire [width_f+3-1:0]fa_fcom,fb_fcom,fs_fcom,fs_fnormalzied;
wire [$clog2(width_total)-1:0]fs_fshiftnumber;

//swap
assign fb_math = {op^fb[31],fb[30:0]};
assign {fa_s,fa_e,fa_f} = (fa[30:23] > fb[30:23])? fa:fb_math;
assign {fb_s,fb_e,fb_f} = (fa[30:23] > fb[30:23])? fb_math:fa;
//extend
assign fa_fex = {3'b001,fa_f};
assign fb_fex = {3'b001,fb_f};
//shift
assign ex_diff = fa_e - fb_e;
assign fb_fexshift = fb_fex >> ex_diff;
//complement
assign fa_fcom = (fa_s)? ~fa_fex+26'd1:fa_fex;
assign fb_fcom = (fb_s)? ~fb_fexshift+26'd1:fb_fexshift;
//adder
assign fs_fcal = fa_fcom + fb_fcom;
//complement get abs value
assign fs_fcom = (fs_fcal[25])? ~fs_fcal+26'd1:fs_fcal;
//normalize
pen32(.din({8'd0,fs_fcom[23:0]}),.dout(fs_fshiftnumber),.valid(valid));
assign fs_s = fs_fcal[25];
assign fs_e = (fs_fcom[24])? fa_e+8'd1:fa_e-(5'd23-fs_fshiftnumber);
assign fs_fnormalzied = fs_fcom << (5'd23-fs_fshiftnumber);
assign fs_f = (fs_fcom[24])? fs_fcom[23:1]:fs_fnormalzied[22:0];
assign zero = (~valid & ~fs_fcom[25] & ~fs_fcom[24]);
assign fs = (zero)? 32'd0:{fs_s,fs_e,fs_f};

endmodule



