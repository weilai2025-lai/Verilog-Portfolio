library verilog;
use verilog.vl_types.all;
entity div_decoder_vlg_check_tst is
    port(
        dout            : in     vl_logic_vector(31 downto 0);
        sampler_rx      : in     vl_logic
    );
end div_decoder_vlg_check_tst;
