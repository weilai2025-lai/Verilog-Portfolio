library verilog;
use verilog.vl_types.all;
entity bounce_avoid_vlg_check_tst is
    port(
        dout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end bounce_avoid_vlg_check_tst;
