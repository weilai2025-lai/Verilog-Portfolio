library verilog;
use verilog.vl_types.all;
entity pencoder_32bit_vlg_vec_tst is
end pencoder_32bit_vlg_vec_tst;
