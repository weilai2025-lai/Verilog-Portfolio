module ffulladd8bit(cin, a, b, s, cout);

input [7:0]a, b;
input cin;
output [7:0]s;
output cout;

wire c;

ffulladd f0(.cin(cin),.a(a[3:0]),.b(b[3:0]),.s(s[3:0]),.cout(c));
ffulladd f1(.cin(c),.a(a[7:4]),.b(b[7:4]),.s(s[7:4]),.cout(cout));

endmodule

