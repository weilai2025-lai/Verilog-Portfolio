library verilog;
use verilog.vl_types.all;
entity D_FF32bit_vlg_sample_tst is
    port(
        clk             : in     vl_logic;
        din             : in     vl_logic_vector(31 downto 0);
        en              : in     vl_logic;
        rst             : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end D_FF32bit_vlg_sample_tst;
