library verilog;
use verilog.vl_types.all;
entity ffulladd8bit_vlg_vec_tst is
end ffulladd8bit_vlg_vec_tst;
