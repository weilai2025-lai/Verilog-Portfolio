library verilog;
use verilog.vl_types.all;
entity Dff_behavioral_vlg_check_tst is
    port(
        q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Dff_behavioral_vlg_check_tst;
