library verilog;
use verilog.vl_types.all;
entity Freq_div_vlg_vec_tst is
end Freq_div_vlg_vec_tst;
