library verilog;
use verilog.vl_types.all;
entity pen32_vlg_vec_tst is
end pen32_vlg_vec_tst;
