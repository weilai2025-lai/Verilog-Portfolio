library verilog;
use verilog.vl_types.all;
entity div_dec_vlg_vec_tst is
end div_dec_vlg_vec_tst;
