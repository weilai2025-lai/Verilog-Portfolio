library verilog;
use verilog.vl_types.all;
entity mux4to1_vlg_check_tst is
    port(
        dout            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux4to1_vlg_check_tst;
