module mux4to1(din, sel, dout);

input [3:0]din;
input [1:0]sel;
output dout;

wire m0_out, m1out;

mux2to1 m0(.a(din[3]),
           .b(din[2]),
			  .sel(sel[0]),
			  .c(m0_out));

mux2to1 m1(.a(din[1]),
           .b(din[0]),
			  .sel(sel[0]),
			  .c(m1_out));

mux2to1 m2(.a(m0_out),
           .b(m1_out),
			  .sel(sel[1]),
			  .c(dout));
endmodule
