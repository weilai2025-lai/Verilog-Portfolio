module mux8to1(din, sel, dout);

input [7:0]din;
input [2:0]sel;

output dout;

wire m0_out, m1_out;

//--我想要自定義腳位,所以先註解掉--
//mux4to1 m0(.din(din[3:0]),
//			  .sel(sel[1:0]),
//			  .dout(m0_out));
//
//mux4to1 m1(.din(din[7:4]),
//			  .sel(sel[1:0]),
//			  .dout(m1_out));
//			  
//mux2to1 m2(.a(m0_out),
//           .b(m1_out),
//			  .sel(sel[2]),
//			  .c(dout));

mux4to1 m0(.din({din[7], din[6], din[5], din[4]}),
           .sel({sel[1], sel[0]}),
			  .dout(m0_out));
			  
mux4to1 m1(.din({din[3], din[2], din[1], din[0]}),
           .sel({sel[1], sel[0]}),
			  .dout(m1_out));
			  
mux2to1 m2(.a(m0_out),
           .b(m1_out),
			  .sel(sel[2]),
			  .c(dout));
			  
endmodule
