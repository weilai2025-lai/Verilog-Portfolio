library verilog;
use verilog.vl_types.all;
entity acc32_vlg_vec_tst is
end acc32_vlg_vec_tst;
