module pen32(din,dout,valid);
parameter width_in = 32;
parameter width_out = 5;

input [width_in-1:0]din;
output reg[width_out-1:0]dout;
output reg valid;
integer i;

always @(*)
begin
	valid = 0;
	dout = 'd0;
	for(i=0;i<32;i=i+1) begin
		if(din[i]) begin
			dout = i;
			valid = 1;
		end
	end
end
endmodule

