library verilog;
use verilog.vl_types.all;
entity PISPO_vlg_vec_tst is
end PISPO_vlg_vec_tst;
