library verilog;
use verilog.vl_types.all;
entity Accumulator_vlg_vec_tst is
end Accumulator_vlg_vec_tst;
