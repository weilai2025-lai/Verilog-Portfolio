library verilog;
use verilog.vl_types.all;
entity D_FF32bit_vlg_vec_tst is
end D_FF32bit_vlg_vec_tst;
