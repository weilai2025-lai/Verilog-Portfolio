library verilog;
use verilog.vl_types.all;
entity D_ff_vlg_vec_tst is
end D_ff_vlg_vec_tst;
