library verilog;
use verilog.vl_types.all;
entity D_Latchbev_vlg_vec_tst is
end D_Latchbev_vlg_vec_tst;
