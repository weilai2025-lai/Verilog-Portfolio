library verilog;
use verilog.vl_types.all;
entity accum_vlg_vec_tst is
end accum_vlg_vec_tst;
