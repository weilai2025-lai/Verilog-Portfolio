library verilog;
use verilog.vl_types.all;
entity count111_mealy_vlg_vec_tst is
end count111_mealy_vlg_vec_tst;
